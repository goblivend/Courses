-- Squelette pour l'exercice RamChip

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity RamChip_tb is
  
end entity;

architecture Bench of RamChip_tb is
   
begin
  

end architecture;
